//
// Gate XOR combinacional
//
module gxor(input a, input b, output y);
  
  assign y = a ^ b;

endmodule

